`define DATA_WIDTH 8
`define CMD_WIDTH  4 
`define no_of_items 20
parameter RESULT_WIDTH = `DATA_WIDTH + 1 ;
