interface alu_assertions(clk,rst,ce,opa,opb,mode,inp_valid,cmd,cin,res,err,cout,oflow,g,l,e);
	input clk;
	input rst;
	input ce;
	input [`DATA_WIDTH - 1 : 0] opa;
	input [`DATA_WIDTH - 1 : 0]opb;
	input mode;
	input [1:0] inp_valid;
	input [`CMD_WIDTH - 1 : 0]cmd;
	input cin;
	input [RESULT_WIDTH - 1 : 0]res;
	input err,cout,oflow,g,l,e;

	property ALU_Known;
		@(posedge clk)
		##1 !($isunknown({rst,ce,opa,opb,mode,inp_valid,cmd,cin}));
	endproperty

	ALU_KNOWN: assert property(ALU_Known)
	$info("INPUTS SIGNALS ARE KNOWN");
	else $info("INPUTS SIGNALS ARE UNKNOWN %d %d %d %d %d %d %d %d",rst,ce,opa,opb,mode,inp_valid,cmd,cin);

	ALU_RESET: assert property(@(posedge clk) ##10 rst )
	$info("RESET IS TRIGGERED");
	else $info("RESET IS NOT TRIGGERED");

	property ALU_Clock_Enable;
		@(posedge clk)
		 !ce |=> ($stable(res));
	endproperty

	ALU_CLOCK_ENABLE: assert property(ALU_Clock_Enable)
  $info("OUTPUTS ARE  LATCHED ");
	else $info("OUTPUTS ARE NOT  LATCHED :%b %d %d %d %d %d %d",res,oflow,cout,g,l,e,err);
endinterface
