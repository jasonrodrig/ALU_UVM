`define DATA_WIDTH 8
`define CMD_WIDTH  4 
`define no_of_items 200 
`define DW 8
`define CW 4
parameter RESULT_WIDTH = `DATA_WIDTH + 1 ;
