alsjdj
